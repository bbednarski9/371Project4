// nios_system.v

<<<<<<< HEAD
// Generated using ACDS version 14.0 200 at 2016.02.22.15:45:24
=======
// Generated using ACDS version 14.0 200 at 2016.02.22.20:35:48
>>>>>>> origin/master

`timescale 1 ps / 1 ps
module nios_system (
		input  wire       reset_reset_n,                //                 reset.reset_n
		output wire [7:0] ledr_export,                  //                  ledr.export
		input  wire [7:0] paralleltoprocessor_export,   //   paralleltoprocessor.export
		input  wire       clk_clk,                      //                   clk.clk
		output wire [7:0] parallelfromprocessor_export, // parallelfromprocessor.export
		output wire       transmitenable_export,        //        transmitenable.export
		output wire       charactersent_export,         //         charactersent.export
		output wire       load_export,                  //                  load.export
		input  wire       characterreceived_export      //     characterreceived.export
	);

	wire         cpu_instruction_master_waitrequest;                          // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [13:0] cpu_instruction_master_address;                              // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                 // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                             // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_data_master_waitrequest;                                 // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                   // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [13:0] cpu_data_master_address;                                     // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire         cpu_data_master_write;                                       // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire         cpu_data_master_read;                                        // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                    // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                                 // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire   [3:0] cpu_data_master_byteenable;                                  // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;         // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;           // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;             // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;               // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;            // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;         // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;          // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;                         // mm_interconnect_0:LEDR_s1_writedata -> LEDR:writedata
	wire   [1:0] mm_interconnect_0_ledr_s1_address;                           // mm_interconnect_0:LEDR_s1_address -> LEDR:address
	wire         mm_interconnect_0_ledr_s1_chipselect;                        // mm_interconnect_0:LEDR_s1_chipselect -> LEDR:chipselect
	wire         mm_interconnect_0_ledr_s1_write;                             // mm_interconnect_0:LEDR_s1_write -> LEDR:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;                          // LEDR:readdata -> mm_interconnect_0:LEDR_s1_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire   [1:0] mm_interconnect_0_paralleltoprocessor_s1_address;            // mm_interconnect_0:ParallelToProcessor_s1_address -> ParallelToProcessor:address
	wire  [31:0] mm_interconnect_0_paralleltoprocessor_s1_readdata;           // ParallelToProcessor:readdata -> mm_interconnect_0:ParallelToProcessor_s1_readdata
	wire  [31:0] mm_interconnect_0_parallelfromprocessor_s1_writedata;        // mm_interconnect_0:ParallelFromProcessor_s1_writedata -> ParallelFromProcessor:writedata
	wire   [1:0] mm_interconnect_0_parallelfromprocessor_s1_address;          // mm_interconnect_0:ParallelFromProcessor_s1_address -> ParallelFromProcessor:address
	wire         mm_interconnect_0_parallelfromprocessor_s1_chipselect;       // mm_interconnect_0:ParallelFromProcessor_s1_chipselect -> ParallelFromProcessor:chipselect
	wire         mm_interconnect_0_parallelfromprocessor_s1_write;            // mm_interconnect_0:ParallelFromProcessor_s1_write -> ParallelFromProcessor:write_n
	wire  [31:0] mm_interconnect_0_parallelfromprocessor_s1_readdata;         // ParallelFromProcessor:readdata -> mm_interconnect_0:ParallelFromProcessor_s1_readdata
	wire  [31:0] mm_interconnect_0_transmitenable_s1_writedata;               // mm_interconnect_0:TransmitEnable_s1_writedata -> TransmitEnable:writedata
	wire   [1:0] mm_interconnect_0_transmitenable_s1_address;                 // mm_interconnect_0:TransmitEnable_s1_address -> TransmitEnable:address
	wire         mm_interconnect_0_transmitenable_s1_chipselect;              // mm_interconnect_0:TransmitEnable_s1_chipselect -> TransmitEnable:chipselect
	wire         mm_interconnect_0_transmitenable_s1_write;                   // mm_interconnect_0:TransmitEnable_s1_write -> TransmitEnable:write_n
	wire  [31:0] mm_interconnect_0_transmitenable_s1_readdata;                // TransmitEnable:readdata -> mm_interconnect_0:TransmitEnable_s1_readdata
	wire  [31:0] mm_interconnect_0_charactersent_s1_writedata;                // mm_interconnect_0:CharacterSent_s1_writedata -> CharacterSent:writedata
	wire   [1:0] mm_interconnect_0_charactersent_s1_address;                  // mm_interconnect_0:CharacterSent_s1_address -> CharacterSent:address
	wire         mm_interconnect_0_charactersent_s1_chipselect;               // mm_interconnect_0:CharacterSent_s1_chipselect -> CharacterSent:chipselect
	wire         mm_interconnect_0_charactersent_s1_write;                    // mm_interconnect_0:CharacterSent_s1_write -> CharacterSent:write_n
	wire  [31:0] mm_interconnect_0_charactersent_s1_readdata;                 // CharacterSent:readdata -> mm_interconnect_0:CharacterSent_s1_readdata
	wire  [31:0] mm_interconnect_0_load_s1_writedata;                         // mm_interconnect_0:Load_s1_writedata -> Load:writedata
	wire   [1:0] mm_interconnect_0_load_s1_address;                           // mm_interconnect_0:Load_s1_address -> Load:address
	wire         mm_interconnect_0_load_s1_chipselect;                        // mm_interconnect_0:Load_s1_chipselect -> Load:chipselect
	wire         mm_interconnect_0_load_s1_write;                             // mm_interconnect_0:Load_s1_write -> Load:write_n
	wire  [31:0] mm_interconnect_0_load_s1_readdata;                          // Load:readdata -> mm_interconnect_0:Load_s1_readdata
	wire   [1:0] mm_interconnect_0_characterreceived_s1_address;              // mm_interconnect_0:CharacterReceived_s1_address -> CharacterReceived:address
	wire  [31:0] mm_interconnect_0_characterreceived_s1_readdata;             // CharacterReceived:readdata -> mm_interconnect_0:CharacterReceived_s1_readdata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] cpu_d_irq_irq;                                               // irq_mapper:sender_irq -> cpu:d_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [CharacterReceived:reset_n, CharacterSent:reset_n, LEDR:reset_n, Load:reset_n, ParallelFromProcessor:reset_n, ParallelToProcessor:reset_n, TransmitEnable:reset_n, cpu:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [cpu:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                           // cpu:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	nios_system_cpu cpu (
		.clk                                   (clk_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	nios_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	nios_system_LEDR ledr (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (ledr_export)                           // external_connection.export
	);

	nios_system_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_system_ParallelToProcessor paralleltoprocessor (
		.clk      (clk_clk),                                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address  (mm_interconnect_0_paralleltoprocessor_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_paralleltoprocessor_s1_readdata), //                    .readdata
		.in_port  (paralleltoprocessor_export)                         // external_connection.export
	);

	nios_system_LEDR parallelfromprocessor (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address    (mm_interconnect_0_parallelfromprocessor_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_parallelfromprocessor_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_parallelfromprocessor_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_parallelfromprocessor_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_parallelfromprocessor_s1_readdata),   //                    .readdata
		.out_port   (parallelfromprocessor_export)                           // external_connection.export
	);

	nios_system_TransmitEnable transmitenable (
		.clk        (clk_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_transmitenable_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_transmitenable_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_transmitenable_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_transmitenable_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_transmitenable_s1_readdata),   //                    .readdata
		.out_port   (transmitenable_export)                           // external_connection.export
	);

	nios_system_TransmitEnable charactersent (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_charactersent_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_charactersent_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_charactersent_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_charactersent_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_charactersent_s1_readdata),   //                    .readdata
		.out_port   (charactersent_export)                           // external_connection.export
	);

	nios_system_TransmitEnable load (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_load_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_load_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_load_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_load_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_load_s1_readdata),   //                    .readdata
		.out_port   (load_export)                           // external_connection.export
	);

	nios_system_CharacterReceived characterreceived (
		.clk      (clk_clk),                                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address  (mm_interconnect_0_characterreceived_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_characterreceived_s1_readdata), //                    .readdata
		.in_port  (characterreceived_export)                         // external_connection.export
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                             (clk_clk),                                                     //                         clk_0_clk.clk
		.cpu_reset_n_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                              // cpu_reset_n_reset_bridge_in_reset.reset
		.cpu_data_master_address                   (cpu_data_master_address),                                     //                   cpu_data_master.address
		.cpu_data_master_waitrequest               (cpu_data_master_waitrequest),                                 //                                  .waitrequest
		.cpu_data_master_byteenable                (cpu_data_master_byteenable),                                  //                                  .byteenable
		.cpu_data_master_read                      (cpu_data_master_read),                                        //                                  .read
		.cpu_data_master_readdata                  (cpu_data_master_readdata),                                    //                                  .readdata
		.cpu_data_master_write                     (cpu_data_master_write),                                       //                                  .write
		.cpu_data_master_writedata                 (cpu_data_master_writedata),                                   //                                  .writedata
		.cpu_data_master_debugaccess               (cpu_data_master_debugaccess),                                 //                                  .debugaccess
		.cpu_instruction_master_address            (cpu_instruction_master_address),                              //            cpu_instruction_master.address
		.cpu_instruction_master_waitrequest        (cpu_instruction_master_waitrequest),                          //                                  .waitrequest
		.cpu_instruction_master_read               (cpu_instruction_master_read),                                 //                                  .read
		.cpu_instruction_master_readdata           (cpu_instruction_master_readdata),                             //                                  .readdata
		.CharacterReceived_s1_address              (mm_interconnect_0_characterreceived_s1_address),              //              CharacterReceived_s1.address
		.CharacterReceived_s1_readdata             (mm_interconnect_0_characterreceived_s1_readdata),             //                                  .readdata
		.CharacterSent_s1_address                  (mm_interconnect_0_charactersent_s1_address),                  //                  CharacterSent_s1.address
		.CharacterSent_s1_write                    (mm_interconnect_0_charactersent_s1_write),                    //                                  .write
		.CharacterSent_s1_readdata                 (mm_interconnect_0_charactersent_s1_readdata),                 //                                  .readdata
		.CharacterSent_s1_writedata                (mm_interconnect_0_charactersent_s1_writedata),                //                                  .writedata
		.CharacterSent_s1_chipselect               (mm_interconnect_0_charactersent_s1_chipselect),               //                                  .chipselect
		.cpu_jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),             //             cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),               //                                  .write
		.cpu_jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),                //                                  .read
		.cpu_jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),            //                                  .readdata
		.cpu_jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),           //                                  .writedata
		.cpu_jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),          //                                  .byteenable
		.cpu_jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),         //                                  .waitrequest
		.cpu_jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),         //                                  .debugaccess
		.jtag_uart_0_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //     jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                  .write
		.jtag_uart_0_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                  .read
		.jtag_uart_0_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                  .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                  .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                  .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                  .chipselect
		.LEDR_s1_address                           (mm_interconnect_0_ledr_s1_address),                           //                           LEDR_s1.address
		.LEDR_s1_write                             (mm_interconnect_0_ledr_s1_write),                             //                                  .write
		.LEDR_s1_readdata                          (mm_interconnect_0_ledr_s1_readdata),                          //                                  .readdata
		.LEDR_s1_writedata                         (mm_interconnect_0_ledr_s1_writedata),                         //                                  .writedata
		.LEDR_s1_chipselect                        (mm_interconnect_0_ledr_s1_chipselect),                        //                                  .chipselect
		.Load_s1_address                           (mm_interconnect_0_load_s1_address),                           //                           Load_s1.address
		.Load_s1_write                             (mm_interconnect_0_load_s1_write),                             //                                  .write
		.Load_s1_readdata                          (mm_interconnect_0_load_s1_readdata),                          //                                  .readdata
		.Load_s1_writedata                         (mm_interconnect_0_load_s1_writedata),                         //                                  .writedata
		.Load_s1_chipselect                        (mm_interconnect_0_load_s1_chipselect),                        //                                  .chipselect
		.onchip_memory2_0_s1_address               (mm_interconnect_0_onchip_memory2_0_s1_address),               //               onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                 (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                  .write
		.onchip_memory2_0_s1_readdata              (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                  .readdata
		.onchip_memory2_0_s1_writedata             (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                  .writedata
		.onchip_memory2_0_s1_byteenable            (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                  .byteenable
		.onchip_memory2_0_s1_chipselect            (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                  .chipselect
		.onchip_memory2_0_s1_clken                 (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                  .clken
		.ParallelFromProcessor_s1_address          (mm_interconnect_0_parallelfromprocessor_s1_address),          //          ParallelFromProcessor_s1.address
		.ParallelFromProcessor_s1_write            (mm_interconnect_0_parallelfromprocessor_s1_write),            //                                  .write
		.ParallelFromProcessor_s1_readdata         (mm_interconnect_0_parallelfromprocessor_s1_readdata),         //                                  .readdata
		.ParallelFromProcessor_s1_writedata        (mm_interconnect_0_parallelfromprocessor_s1_writedata),        //                                  .writedata
		.ParallelFromProcessor_s1_chipselect       (mm_interconnect_0_parallelfromprocessor_s1_chipselect),       //                                  .chipselect
		.ParallelToProcessor_s1_address            (mm_interconnect_0_paralleltoprocessor_s1_address),            //            ParallelToProcessor_s1.address
		.ParallelToProcessor_s1_readdata           (mm_interconnect_0_paralleltoprocessor_s1_readdata),           //                                  .readdata
		.TransmitEnable_s1_address                 (mm_interconnect_0_transmitenable_s1_address),                 //                 TransmitEnable_s1.address
		.TransmitEnable_s1_write                   (mm_interconnect_0_transmitenable_s1_write),                   //                                  .write
		.TransmitEnable_s1_readdata                (mm_interconnect_0_transmitenable_s1_readdata),                //                                  .readdata
		.TransmitEnable_s1_writedata               (mm_interconnect_0_transmitenable_s1_writedata),               //                                  .writedata
		.TransmitEnable_s1_chipselect              (mm_interconnect_0_transmitenable_s1_chipselect)               //                                  .chipselect
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
