
module nios_system (
	reset_reset_n,
	ledr_export,
	clk_clk);	

	input		reset_reset_n;
	output	[7:0]	ledr_export;
	input		clk_clk;
endmodule
